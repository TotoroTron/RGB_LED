library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package parameters is
    type table is array(0 to 63) of integer;
    type table255 is array(0 to 255) of integer;
    signal gamma : table :=
    (
        0, 0, 0, 0, 0, 0, 0, 1,
        1, 1, 1, 1, 2, 2, 2, 3, 
        3, 4, 4, 5, 5, 6, 6, 7,
        8, 8, 9, 10, 11, 11, 12, 13,
        14, 15, 16, 17, 18, 20, 21, 22,
        23, 24, 26, 27, 29, 30, 32, 33, 
        35, 36, 38, 40, 41, 43, 45, 47, 
        49, 51, 53, 55, 57, 59, 61, 63
    );
    
    signal gamma255 : table255 :=
    (
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
        0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1,
        1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2,
        2, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 5, 5, 5,
        5, 6, 6, 6, 6, 7, 7, 7, 7, 8, 8, 8, 9, 9, 9, 10,
        10, 10, 11, 11, 11, 12, 12, 13, 13, 13, 14, 14, 15, 15, 16, 16,
        17, 17, 18, 18, 19, 19, 20, 20, 21, 21, 22, 22, 23, 24, 24, 25,
        25, 26, 27, 27, 28, 29, 29, 30, 31, 32, 32, 33, 34, 35, 35, 36,
        37, 38, 39, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 50,
        51, 52, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 66, 67, 68,
        69, 70, 72, 73, 74, 75, 77, 78, 79, 81, 82, 83, 85, 86, 87, 89,
        90, 92, 93, 95, 96, 98, 99,101,102,104,105,107,109,110,112,114,
        115,117,119,120,122,124,126,127,129,131,133,135,137,138,140,142,
        144,146,148,150,152,154,156,158,160,162,164,167,169,171,173,175,
        177,180,182,184,186,189,191,193,196,198,200,203,205,208,210,213,
        215,218,220,223,225,228,231,233,236,239,241,244,247,249,252,255
    );
    
    constant IMG_WIDTH : integer := 32;
    constant IMG_HEIGHT : integer := 32;
    constant COLOR_DEPTH : integer := 24;
    constant NUM_FRAMES : integer := 29;
    constant IMG_FILE : string := "rainbow2.mem";

end package;
